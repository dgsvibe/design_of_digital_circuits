library verilog;
use verilog.vl_types.all;
entity pnand_vlg_vec_tst is
end pnand_vlg_vec_tst;
