library verilog;
use verilog.vl_types.all;
entity reg10b_vlg_check_tst is
    port(
        q               : in     vl_logic_vector(9 downto 0);
        sampler_rx      : in     vl_logic
    );
end reg10b_vlg_check_tst;
