LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mux_2x1 IS
PORT(	e0, e1: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		sel: IN STD_LOGIC;
		s: OUT STD_LOGIC_VECTOR(9 DOWNTO 0));
END mux_2x1;

ARCHITECTURE behavioral OF mux_2x1 IS
BEGIN
s <= e0 WHEN (sel = '0') ELSE e1;
END behavioral;