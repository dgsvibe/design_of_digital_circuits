library verilog;
use verilog.vl_types.all;
entity dbreg_vlg_vec_tst is
end dbreg_vlg_vec_tst;
