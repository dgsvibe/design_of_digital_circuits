library verilog;
use verilog.vl_types.all;
entity reg10bhlb_vlg_vec_tst is
end reg10bhlb_vlg_vec_tst;
