library verilog;
use verilog.vl_types.all;
entity reg10b_vlg_vec_tst is
end reg10b_vlg_vec_tst;
