library verilog;
use verilog.vl_types.all;
entity Sub1_structural_vlg_check_tst is
    port(
        S               : in     vl_logic_vector(9 downto 0);
        sampler_rx      : in     vl_logic
    );
end Sub1_structural_vlg_check_tst;
