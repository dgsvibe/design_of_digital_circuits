library verilog;
use verilog.vl_types.all;
entity pnand_vlg_check_tst is
    port(
        s               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end pnand_vlg_check_tst;
