library verilog;
use verilog.vl_types.all;
entity pnot_vlg_vec_tst is
end pnot_vlg_vec_tst;
