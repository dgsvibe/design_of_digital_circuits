library verilog;
use verilog.vl_types.all;
entity Sub1_structural_vlg_vec_tst is
end Sub1_structural_vlg_vec_tst;
