library verilog;
use verilog.vl_types.all;
entity exercicio01 is
    port(
        s9              : out    vl_logic;
        rst             : in     vl_logic;
        ck              : in     vl_logic;
        c9              : in     vl_logic;
        c0              : in     vl_logic;
        c1              : in     vl_logic;
        c2              : in     vl_logic;
        c3              : in     vl_logic;
        c4              : in     vl_logic;
        c5              : in     vl_logic;
        c6              : in     vl_logic;
        c7              : in     vl_logic;
        c8              : in     vl_logic;
        s8              : out    vl_logic;
        s7              : out    vl_logic;
        s6              : out    vl_logic;
        s5              : out    vl_logic;
        s4              : out    vl_logic;
        s3              : out    vl_logic;
        s2              : out    vl_logic;
        s1              : out    vl_logic;
        s0              : out    vl_logic
    );
end exercicio01;
