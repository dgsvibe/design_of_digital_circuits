library verilog;
use verilog.vl_types.all;
entity Sub1_behavioral_vlg_vec_tst is
end Sub1_behavioral_vlg_vec_tst;
