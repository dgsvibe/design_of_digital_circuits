LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY e2mod IS
PORT(	enter: IN STD_LOGIC;
		data: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		s: OUT STD_LOGIC_VECTOR(9 DOWNTO 0));
END e2mod;

ARCHITECTURE arch OF e2mod IS
BEGIN
	p: PROCESS(enter, data) BEGIN
		IF(enter='1') THEN s(9 DOWNTO 0)<=data(9 DOWNTO 0); 
		END IF;
	END PROCESS p;
END arch;