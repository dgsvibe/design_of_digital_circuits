library verilog;
use verilog.vl_types.all;
entity exercicio01_vlg_sample_tst is
    port(
        c0              : in     vl_logic;
        c1              : in     vl_logic;
        c2              : in     vl_logic;
        c3              : in     vl_logic;
        c4              : in     vl_logic;
        c5              : in     vl_logic;
        c6              : in     vl_logic;
        c7              : in     vl_logic;
        c8              : in     vl_logic;
        c9              : in     vl_logic;
        ck              : in     vl_logic;
        rst             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end exercicio01_vlg_sample_tst;
