library verilog;
use verilog.vl_types.all;
entity mtfffixed_vlg_vec_tst is
end mtfffixed_vlg_vec_tst;
