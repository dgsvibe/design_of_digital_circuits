library verilog;
use verilog.vl_types.all;
entity exercicio01_vlg_vec_tst is
end exercicio01_vlg_vec_tst;
