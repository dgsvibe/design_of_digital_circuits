library verilog;
use verilog.vl_types.all;
entity demux2x1_vlg_vec_tst is
end demux2x1_vlg_vec_tst;
