LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY pnot IS
PORT(	a: IN STD_LOGIC;
		s: OUT STD_LOGIC);
END pnot;

ARCHITECTURE arch OF pnot IS
BEGIN
s<=NOT(a);
END arch;