library verilog;
use verilog.vl_types.all;
entity dff_behavioral_vlg_check_tst is
    port(
        q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end dff_behavioral_vlg_check_tst;
