LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY Mux2x1x10 IS
	PORT(	e0: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
			e1: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
			c: IN STD_LOGIC;
			s: OUT STD_LOGIC_VECTOR(9 DOWNTO 0));
END Mux2x1x10;

ARCHITECTURE arch OF Mux2x1x10 IS
BEGIN
	p: PROCESS(e0, e1, c)
	BEGIN
		IF(c='0') THEN s(9 DOWNTO 0)<=e0(9 DOWNTO 0);
			ELSIF(c='1') THEN s(9 DOWNTO 0)<=e1(9 DOWNTO 0);
		END IF;
	END PROCESS;
	
END arch;