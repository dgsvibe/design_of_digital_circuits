library verilog;
use verilog.vl_types.all;
entity reg6b_vlg_vec_tst is
end reg6b_vlg_vec_tst;
