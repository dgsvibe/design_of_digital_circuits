library verilog;
use verilog.vl_types.all;
entity Mux2x1x6_vlg_vec_tst is
end Mux2x1x6_vlg_vec_tst;
