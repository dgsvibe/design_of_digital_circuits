library verilog;
use verilog.vl_types.all;
entity exercicio02_vlg_vec_tst is
end exercicio02_vlg_vec_tst;
