library verilog;
use verilog.vl_types.all;
entity e2mod_vlg_vec_tst is
end e2mod_vlg_vec_tst;
