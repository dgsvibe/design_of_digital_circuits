library verilog;
use verilog.vl_types.all;
entity sum6b_vlg_vec_tst is
end sum6b_vlg_vec_tst;
