library verilog;
use verilog.vl_types.all;
entity flipflopt_vlg_vec_tst is
end flipflopt_vlg_vec_tst;
