library verilog;
use verilog.vl_types.all;
entity exercicio01_vlg_check_tst is
    port(
        s0              : in     vl_logic;
        s1              : in     vl_logic;
        s2              : in     vl_logic;
        s3              : in     vl_logic;
        s4              : in     vl_logic;
        s5              : in     vl_logic;
        s6              : in     vl_logic;
        s7              : in     vl_logic;
        s8              : in     vl_logic;
        s9              : in     vl_logic;
        sginal_nor      : in     vl_logic;
        signal_T        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end exercicio01_vlg_check_tst;
