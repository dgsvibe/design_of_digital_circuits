library verilog;
use verilog.vl_types.all;
entity sum10b_vlg_vec_tst is
end sum10b_vlg_vec_tst;
