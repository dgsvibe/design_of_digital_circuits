library verilog;
use verilog.vl_types.all;
entity dff_behavioral_vlg_vec_tst is
end dff_behavioral_vlg_vec_tst;
